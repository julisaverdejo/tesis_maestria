// Author: Julisa Verdejo Palacios
// Name: rom_volts.v
//
// Description: 


module rom_volts (
  input      [4:0] addr_i,
  output reg [11:0] rom_o
);

  always@(addr_i)  
    case(addr_i)
       0 : rom_o = 12'b000000000000; //0.00
       1 : rom_o = 12'b000001111100; //0.10
       2 : rom_o = 12'b000011111000; //0.20
       3 : rom_o = 12'b000101110100; //0.30
       4 : rom_o = 12'b000111110000; //0.40
       5 : rom_o = 12'b001001101100; //0.50
       6 : rom_o = 12'b001011101000; //0.60
       7 : rom_o = 12'b001101100100; //0.70
       8 : rom_o = 12'b001111100000; //0.80
       9 : rom_o = 12'b010001011100; //0.90
      10 : rom_o = 12'b010011011000; //1.00
      11 : rom_o = 12'b010101010100; //1.10
      12 : rom_o = 12'b010111010000; //1.20
      13 : rom_o = 12'b011001001100; //1.30
      14 : rom_o = 12'b011011001000; //1.40
      15 : rom_o = 12'b011101000100; //1.50
      16 : rom_o = 12'b011111000000; //1.60
      17 : rom_o = 12'b100000111100; //1.70
      18 : rom_o = 12'b100010111000; //1.80
      19 : rom_o = 12'b100100110100; //1.90
      20 : rom_o = 12'b100110110000; //2.00
      21 : rom_o = 12'b101000101100; //2.10
      22 : rom_o = 12'b101010101000; //2.20
      23 : rom_o = 12'b101100100100; //2.30
      24 : rom_o = 12'b101110100000; //2.40
      25 : rom_o = 12'b110000011100; //2.50
      26 : rom_o = 12'b110010011000; //2.60
      27 : rom_o = 12'b110100010100; //2.70
      28 : rom_o = 12'b110110010000; //2.80
      29 : rom_o = 12'b111000001100; //2.90
      30 : rom_o = 12'b111010001000; //3.00	  
	  default: rom_o = 12'b000000000000;
	endcase
endmodule